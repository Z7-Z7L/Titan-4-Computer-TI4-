module IO (
  
);
  
endmodule