module Mem (
  
);
  
endmodule